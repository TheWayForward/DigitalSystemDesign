//breath_multifunction
module breath_multifunction(
	clk,
	rst,
	led
);

	//basic
	input clk,rst;
	output led;

	
	
endmodule
